`timescale 1 ns / 1 ps

module pixelTop_tb;
   logic clk =0;
   logic reset =0;
   logic start =0;
   parameter integer clk_period = 50;
   parameter integer sim_end = clk_period*2400;
   always #clk_period clk=~clk;

   PIXEL_TOP pixeltop(.clk(clk), .reset(reset), .start(start));

   initial
     begin
        reset = 1;

        #clk_period  reset=0;

        $dumpfile("pixelTop_tb.vcd");
        $dumpvars(0,pixelTop_tb);

        #2000 start = 1;

        #clk_period  start=0;


        #57000 reset = 1;
        #200  reset = 0;

        #1000 start = 1;
        #clk_period  start=0;


        #25000 reset = 1;
        #clk_period  reset=0;



        

        #sim_end
          $stop;
     end

endmodule
